-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Wed May 17 20:31:26 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ControlSystemUnit IS
    PORT (
        reset : IN STD_LOGIC;
        clock : IN STD_LOGIC;
        start : IN STD_LOGIC;
        freezeEnd : IN STD_LOGIC;
        extraEn : IN STD_LOGIC;
        newPrg : IN STD_LOGIC;
        freeze : IN STD_LOGIC;
        en_1 : OUT STD_LOGIC;
        en_2 : OUT STD_LOGIC;
        en_3 : OUT STD_LOGIC;
        start_stop : OUT STD_LOGIC;
        freezeStart : OUT STD_LOGIC;
        rstGlobal : OUT STD_LOGIC
    );
END ControlSystemUnit;

ARCHITECTURE BEHAVIOR OF ControlSystemUnit IS
    TYPE type_fstate IS (Init,Menu,Timer,TimeProcess,StartPrg,Stop,Extra);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN

    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,start,freezeEnd,extraEn,newPrg,freeze)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Init;
            en_1 <= '0';
            en_2 <= '0';
            en_3 <= '0';
            start_stop <= '0';
            freezeStart <= '0';
            rstGlobal <= '0';
        ELSE
            en_1 <= '0';
            en_2 <= '0';
            en_3 <= '0';
            start_stop <= '0';
            freezeStart <= '0';
            rstGlobal <= '0';
				
            CASE fstate IS
                WHEN Init =>
                    reg_fstate <= Menu;

                    en_3 <= '0';

                    en_1 <= '0';

                    rstGlobal <= '1';

                    start_stop <= '0';

                    en_2 <= '0';

                    freezeStart <= '0';
                WHEN Menu =>
                    IF ((freeze = '1')) THEN
                        reg_fstate <= Timer;
                    ELSIF (start = '1') THEN
                        reg_fstate <= StartPrg;
                    ELSE
                        reg_fstate <= Menu;
                    END IF;
                    en_3 <= '0';

                    en_1 <= '1';

                    rstGlobal <= '0';

                    start_stop <= '0';

                    en_2 <= '0';

                    freezeStart <= '0';
						  
                WHEN Timer =>
                    IF (((start = '1') AND NOT((freeze = '1')))) THEN
                        reg_fstate <= TimeProcess;
                    ELSE
                        reg_fstate <= Timer;
                    END IF;

                    en_3 <= '1';

                    en_1 <= '1';

                    rstGlobal <= '0';

                    start_stop <= '0';

                    en_2 <= '0';

                    freezeStart <= '0';
						  
                WHEN TimeProcess =>
					 
                    IF (freezeEnd = '1') THEN
                        reg_fstate <= StartPrg;
                    ELSE
                        reg_fstate <= TimeProcess;
                    END IF;

                    en_3 <= '1';

                    en_1 <= '0';

                    rstGlobal <= '0';

                    start_stop <= '0';

                    en_2 <= '0';

                    freezeStart <= '1';
                WHEN StartPrg =>
                    IF (start = '1') THEN
                        reg_fstate <= Stop;
                    ELSIF (extraEn = '1') THEN
                        reg_fstate <= Extra;
                    ELSIF (newPrg = '1') THEN
                        reg_fstate <= Init;
                    ELSE
                        reg_fstate <= StartPrg;
                    END IF;

                    en_3 <= '0';

                    en_1 <= '0';

                    rstGlobal <= '0';

                    start_stop <= '1';

                    en_2 <= '0';

                    freezeStart <= '0';
                WHEN Stop =>
                    IF (start = '1') THEN
                        reg_fstate <= StartPrg;
                    ELSE
                        reg_fstate <= Stop;
                    END IF;

                    en_3 <= '0';

                    en_1 <= '0';

                    rstGlobal <= '0';

                    en_2 <= '0';

                    freezeStart <= '0';
                WHEN Extra =>
                    IF (start = '1') THEN
                        reg_fstate <= StartPrg;
                    ELSE
                        reg_fstate <= Extra;
                    END IF;

                    en_3 <= '0';

                    en_1 <= '0';

                    rstGlobal <= '0';

                    start_stop <= '0';

                    en_2 <= '1';

                    freezeStart <= '0';
                WHEN OTHERS =>
                    en_1 <= 'X';
                    en_2 <= 'X';
                    en_3 <= 'X';
                    start_stop <= 'X';
                    freezeStart <= 'X';
                    rstGlobal <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
